`define PCKG_SZ 32 
`define DRVRS 4 
`define BITS 1

